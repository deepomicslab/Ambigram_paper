chrom_5p	bkpos_5p	strand_5p	chrom_3p	bkpos_3p	strand_3p	avg_cn
chr7	54605701	+	chr7	55191871	+	30.6096319717
chr7	55201724	+	chr7	55222812	+	28.4734917157
chr7	55191871	+	chr7	55223396	+	23.285007155
chr7	54706322	+	chr7	55201725	+	195.842655989
chr7	55289061	+	chr7	54706322	+	179.298444894